library verilog;
use verilog.vl_types.all;
entity CPUDesign_vlg_vec_tst is
end CPUDesign_vlg_vec_tst;
